magic
tech sky130A
magscale 1 2
timestamp 1707999654
<< metal1 >>
rect 22108 22494 22118 22606
rect 22252 22494 22262 22606
rect 22498 22500 22508 22612
rect 22642 22500 22652 22612
rect 23132 22512 23142 22624
rect 23276 22512 23286 22624
rect 23770 22512 23780 22624
rect 23914 22512 23924 22624
rect 22120 22008 22204 22494
rect 22528 22132 22612 22500
rect 23158 22226 23242 22512
rect 23158 22142 23298 22226
rect 22528 22048 22972 22132
rect 22120 21924 22596 22008
rect 21392 21193 22287 21311
rect 22512 21198 22596 21924
rect 22888 21198 22972 22048
rect 23214 21196 23298 22142
rect 23804 21764 23888 22512
rect 23618 21680 23888 21764
rect 23618 21204 23702 21680
rect 21048 20848 21058 21090
rect 21304 21020 21314 21090
rect 21392 21020 21510 21193
rect 21304 20902 21510 21020
rect 21304 20848 21314 20902
rect 22140 17734 22614 18118
rect 22874 17851 22960 17870
rect 23206 17853 23292 17862
rect 22228 15189 22333 17734
rect 22874 17722 22961 17851
rect 22875 17653 22961 17722
rect 22558 17567 22961 17653
rect 23205 17714 23292 17853
rect 23614 17859 23700 17862
rect 23614 17714 23705 17859
rect 25784 17788 25794 17888
rect 25906 17788 25916 17888
rect 22558 17384 22644 17567
rect 22552 15189 22650 15414
rect 22729 15339 22815 17567
rect 23205 17554 23291 17714
rect 23619 17565 23705 17714
rect 25787 17565 25873 17788
rect 23619 17556 25873 17565
rect 23004 17468 23291 17554
rect 23004 17406 23090 17468
rect 22729 15253 23101 15339
rect 23205 15331 23291 17468
rect 23438 17479 25873 17556
rect 23438 17470 23705 17479
rect 23438 17408 23524 17470
rect 23205 15245 23507 15331
rect 22228 15091 22650 15189
rect 22228 15088 22333 15091
<< via1 >>
rect 22118 22494 22252 22606
rect 22508 22500 22642 22612
rect 23142 22512 23276 22624
rect 23780 22512 23914 22624
rect 21058 20848 21304 21090
rect 25794 17788 25906 17888
<< metal2 >>
rect 23142 22624 23276 22634
rect 22118 22606 22252 22616
rect 22118 22484 22252 22494
rect 22508 22612 22642 22622
rect 23142 22502 23276 22512
rect 23780 22624 23914 22634
rect 23780 22502 23914 22512
rect 22508 22490 22642 22500
rect 21058 21090 21304 21100
rect 21058 20838 21304 20848
rect 25794 17888 25906 17898
rect 25794 17778 25906 17788
<< via2 >>
rect 22118 22494 22252 22606
rect 22508 22500 22642 22612
rect 23142 22512 23276 22624
rect 23780 22512 23914 22624
rect 21058 20848 21304 21090
rect 25794 17788 25906 17888
<< metal3 >>
rect 23132 22624 23286 22629
rect 22498 22612 22652 22617
rect 22108 22606 22262 22611
rect 22108 22494 22118 22606
rect 22252 22494 22262 22606
rect 22498 22500 22508 22612
rect 22642 22500 22652 22612
rect 23132 22512 23142 22624
rect 23276 22512 23286 22624
rect 23132 22507 23286 22512
rect 23770 22624 23924 22629
rect 23770 22512 23780 22624
rect 23914 22512 23924 22624
rect 23770 22507 23924 22512
rect 22498 22495 22652 22500
rect 22108 22489 22262 22494
rect 21048 21090 21314 21095
rect 21048 20848 21058 21090
rect 21304 20848 21314 21090
rect 21048 20843 21314 20848
rect 25784 17888 25916 17893
rect 25784 17788 25794 17888
rect 25906 17788 25916 17888
rect 25784 17783 25916 17788
<< via3 >>
rect 22118 22494 22252 22606
rect 22508 22500 22642 22612
rect 23142 22512 23276 22624
rect 23780 22512 23914 22624
rect 21058 20848 21304 21090
rect 25794 17788 25906 17888
<< metal4 >>
rect 200 200 500 45152
rect 798 44952 858 45152
rect 1534 44952 1594 45152
rect 2270 44952 2330 45152
rect 3006 44952 3066 45152
rect 3742 44952 3802 45152
rect 4478 44952 4538 45152
rect 5214 44952 5274 45152
rect 5950 44952 6010 45152
rect 6686 44952 6746 45152
rect 7422 44952 7482 45152
rect 8158 44952 8218 45152
rect 8894 44952 8954 45152
rect 9630 44952 9690 45152
rect 9800 21112 10100 45152
rect 10366 44952 10426 45152
rect 11102 44952 11162 45152
rect 11838 44952 11898 45152
rect 12574 44952 12634 45152
rect 13310 44952 13370 45152
rect 14046 44952 14106 45152
rect 14782 44952 14842 45152
rect 15518 44952 15578 45152
rect 16254 44952 16314 45152
rect 16990 44952 17050 45152
rect 17726 44952 17786 45152
rect 18462 44952 18522 45152
rect 19198 44952 19258 45152
rect 19934 44952 19994 45152
rect 20670 44952 20730 45152
rect 21406 44952 21466 45152
rect 22142 44952 22202 45152
rect 22878 44952 22938 45152
rect 23614 44952 23674 45152
rect 24350 44952 24410 45152
rect 25086 44952 25146 45152
rect 25822 44952 25882 45152
rect 26558 44952 26618 45152
rect 27294 26762 27354 45152
rect 22150 26702 27354 26762
rect 22150 22607 22210 26702
rect 28030 26092 28090 45152
rect 22550 26032 28090 26092
rect 22550 22613 22610 26032
rect 28766 25374 28826 45152
rect 23182 25314 28826 25374
rect 23182 22625 23242 25314
rect 29502 24882 29562 45152
rect 30238 44952 30298 45152
rect 30974 44952 31034 45152
rect 31710 44952 31770 45152
rect 23814 24822 29562 24882
rect 23814 22625 23874 24822
rect 23141 22624 23277 22625
rect 22507 22612 22643 22613
rect 22117 22606 22253 22607
rect 22117 22494 22118 22606
rect 22252 22494 22253 22606
rect 22507 22500 22508 22612
rect 22642 22500 22643 22612
rect 23141 22512 23142 22624
rect 23276 22512 23277 22624
rect 23141 22511 23277 22512
rect 23779 22624 23915 22625
rect 23779 22512 23780 22624
rect 23914 22512 23915 22624
rect 23779 22511 23915 22512
rect 22507 22499 22643 22500
rect 22117 22493 22253 22494
rect 9800 21090 21332 21112
rect 9800 20848 21058 21090
rect 21304 20848 21332 21090
rect 9800 20812 21332 20848
rect 200 0 520 200
rect 4816 0 4936 200
rect 9232 0 9352 200
rect 9800 0 10100 20812
rect 25775 17888 31435 17903
rect 25775 17788 25794 17888
rect 25906 17788 31435 17888
rect 25775 17777 31435 17788
rect 31309 1653 31435 17777
rect 13648 0 13768 200
rect 18064 0 18184 200
rect 22480 0 22600 200
rect 26896 0 27016 200
rect 31312 0 31432 1653
use sky130_fd_pr__res_generic_po_6GTJ3K  sky130_fd_pr__res_generic_po_6GTJ3K_0
timestamp 1707999010
transform 1 0 22601 0 1 16365
box -33 -1115 33 1115
use sky130_fd_pr__res_generic_po_6GTJ3K  sky130_fd_pr__res_generic_po_6GTJ3K_1
timestamp 1707999010
transform 1 0 23041 0 1 16363
box -33 -1115 33 1115
use sky130_fd_pr__res_generic_po_6GTJ3K  sky130_fd_pr__res_generic_po_6GTJ3K_2
timestamp 1707999010
transform 1 0 23473 0 1 16377
box -33 -1115 33 1115
use sky130_fd_pr__res_generic_po_M7V662  sky130_fd_pr__res_generic_po_M7V662_0
timestamp 1707999010
transform 1 0 22229 0 1 19523
box -33 -1799 33 1799
use sky130_fd_pr__res_generic_po_M7V662  sky130_fd_pr__res_generic_po_M7V662_1
timestamp 1707999010
transform 1 0 22551 0 1 19531
box -33 -1799 33 1799
use sky130_fd_pr__res_generic_po_M7V662  sky130_fd_pr__res_generic_po_M7V662_2
timestamp 1707999010
transform 1 0 22915 0 1 19527
box -33 -1799 33 1799
use sky130_fd_pr__res_generic_po_M7V662  sky130_fd_pr__res_generic_po_M7V662_3
timestamp 1707999010
transform 1 0 23249 0 1 19515
box -33 -1799 33 1799
use sky130_fd_pr__res_generic_po_M7V662  sky130_fd_pr__res_generic_po_M7V662_4
timestamp 1707999010
transform 1 0 23653 0 1 19519
box -33 -1799 33 1799
<< labels >>
flabel metal4 s 30974 44952 31034 45152 0 FreeSans 480 90 0 0 clk
port 0 nsew signal input
flabel metal4 s 31710 44952 31770 45152 0 FreeSans 480 90 0 0 ena
port 1 nsew signal input
flabel metal4 s 30238 44952 30298 45152 0 FreeSans 480 90 0 0 rst_n
port 2 nsew signal input
flabel metal4 s 31312 0 31432 200 0 FreeSans 960 0 0 0 ua[0]
port 3 nsew signal bidirectional
flabel metal4 s 26896 0 27016 200 0 FreeSans 960 0 0 0 ua[1]
port 4 nsew signal bidirectional
flabel metal4 s 22480 0 22600 200 0 FreeSans 960 0 0 0 ua[2]
port 5 nsew signal bidirectional
flabel metal4 s 18064 0 18184 200 0 FreeSans 960 0 0 0 ua[3]
port 6 nsew signal bidirectional
flabel metal4 s 13648 0 13768 200 0 FreeSans 960 0 0 0 ua[4]
port 7 nsew signal bidirectional
flabel metal4 s 9232 0 9352 200 0 FreeSans 960 0 0 0 ua[5]
port 8 nsew signal bidirectional
flabel metal4 s 4816 0 4936 200 0 FreeSans 960 0 0 0 ua[6]
port 9 nsew signal bidirectional
flabel metal4 s 400 0 520 200 0 FreeSans 960 0 0 0 ua[7]
port 10 nsew signal bidirectional
flabel metal4 s 29502 44952 29562 45152 0 FreeSans 480 90 0 0 ui_in[0]
port 11 nsew signal input
flabel metal4 s 28766 44952 28826 45152 0 FreeSans 480 90 0 0 ui_in[1]
port 12 nsew signal input
flabel metal4 s 28030 44952 28090 45152 0 FreeSans 480 90 0 0 ui_in[2]
port 13 nsew signal input
flabel metal4 s 27294 44952 27354 45152 0 FreeSans 480 90 0 0 ui_in[3]
port 14 nsew signal input
flabel metal4 s 26558 44952 26618 45152 0 FreeSans 480 90 0 0 ui_in[4]
port 15 nsew signal input
flabel metal4 s 25822 44952 25882 45152 0 FreeSans 480 90 0 0 ui_in[5]
port 16 nsew signal input
flabel metal4 s 25086 44952 25146 45152 0 FreeSans 480 90 0 0 ui_in[6]
port 17 nsew signal input
flabel metal4 s 24350 44952 24410 45152 0 FreeSans 480 90 0 0 ui_in[7]
port 18 nsew signal input
flabel metal4 s 23614 44952 23674 45152 0 FreeSans 480 90 0 0 uio_in[0]
port 19 nsew signal input
flabel metal4 s 22878 44952 22938 45152 0 FreeSans 480 90 0 0 uio_in[1]
port 20 nsew signal input
flabel metal4 s 22142 44952 22202 45152 0 FreeSans 480 90 0 0 uio_in[2]
port 21 nsew signal input
flabel metal4 s 21406 44952 21466 45152 0 FreeSans 480 90 0 0 uio_in[3]
port 22 nsew signal input
flabel metal4 s 20670 44952 20730 45152 0 FreeSans 480 90 0 0 uio_in[4]
port 23 nsew signal input
flabel metal4 s 19934 44952 19994 45152 0 FreeSans 480 90 0 0 uio_in[5]
port 24 nsew signal input
flabel metal4 s 19198 44952 19258 45152 0 FreeSans 480 90 0 0 uio_in[6]
port 25 nsew signal input
flabel metal4 s 18462 44952 18522 45152 0 FreeSans 480 90 0 0 uio_in[7]
port 26 nsew signal input
flabel metal4 s 5950 44952 6010 45152 0 FreeSans 480 90 0 0 uio_oe[0]
port 27 nsew signal tristate
flabel metal4 s 5214 44952 5274 45152 0 FreeSans 480 90 0 0 uio_oe[1]
port 28 nsew signal tristate
flabel metal4 s 4478 44952 4538 45152 0 FreeSans 480 90 0 0 uio_oe[2]
port 29 nsew signal tristate
flabel metal4 s 3742 44952 3802 45152 0 FreeSans 480 90 0 0 uio_oe[3]
port 30 nsew signal tristate
flabel metal4 s 3006 44952 3066 45152 0 FreeSans 480 90 0 0 uio_oe[4]
port 31 nsew signal tristate
flabel metal4 s 2270 44952 2330 45152 0 FreeSans 480 90 0 0 uio_oe[5]
port 32 nsew signal tristate
flabel metal4 s 1534 44952 1594 45152 0 FreeSans 480 90 0 0 uio_oe[6]
port 33 nsew signal tristate
flabel metal4 s 798 44952 858 45152 0 FreeSans 480 90 0 0 uio_oe[7]
port 34 nsew signal tristate
flabel metal4 s 11838 44952 11898 45152 0 FreeSans 480 90 0 0 uio_out[0]
port 35 nsew signal tristate
flabel metal4 s 11102 44952 11162 45152 0 FreeSans 480 90 0 0 uio_out[1]
port 36 nsew signal tristate
flabel metal4 s 10366 44952 10426 45152 0 FreeSans 480 90 0 0 uio_out[2]
port 37 nsew signal tristate
flabel metal4 s 9630 44952 9690 45152 0 FreeSans 480 90 0 0 uio_out[3]
port 38 nsew signal tristate
flabel metal4 s 8894 44952 8954 45152 0 FreeSans 480 90 0 0 uio_out[4]
port 39 nsew signal tristate
flabel metal4 s 8158 44952 8218 45152 0 FreeSans 480 90 0 0 uio_out[5]
port 40 nsew signal tristate
flabel metal4 s 7422 44952 7482 45152 0 FreeSans 480 90 0 0 uio_out[6]
port 41 nsew signal tristate
flabel metal4 s 6686 44952 6746 45152 0 FreeSans 480 90 0 0 uio_out[7]
port 42 nsew signal tristate
flabel metal4 s 17726 44952 17786 45152 0 FreeSans 480 90 0 0 uo_out[0]
port 43 nsew signal tristate
flabel metal4 s 16990 44952 17050 45152 0 FreeSans 480 90 0 0 uo_out[1]
port 44 nsew signal tristate
flabel metal4 s 16254 44952 16314 45152 0 FreeSans 480 90 0 0 uo_out[2]
port 45 nsew signal tristate
flabel metal4 s 15518 44952 15578 45152 0 FreeSans 480 90 0 0 uo_out[3]
port 46 nsew signal tristate
flabel metal4 s 14782 44952 14842 45152 0 FreeSans 480 90 0 0 uo_out[4]
port 47 nsew signal tristate
flabel metal4 s 14046 44952 14106 45152 0 FreeSans 480 90 0 0 uo_out[5]
port 48 nsew signal tristate
flabel metal4 s 13310 44952 13370 45152 0 FreeSans 480 90 0 0 uo_out[6]
port 49 nsew signal tristate
flabel metal4 s 12574 44952 12634 45152 0 FreeSans 480 90 0 0 uo_out[7]
port 50 nsew signal tristate
flabel metal4 200 0 500 45152 1 FreeSans 2 0 0 0 VPWR
port 51 nsew power bidirectional
flabel metal4 9800 0 10100 45152 1 FreeSans 2 0 0 0 VGND
port 52 nsew ground bidirectional
<< properties >>
string FIXED_BBOX 0 0 32200 45152
<< end >>
